module test_x(output b);
    assign b = 1'bx;
endmodule

module test_z(output b);
    assign b = 1'bz;
endmodule